module ALU_Control
(
    input wire [1:0] alu_op,
    input wire [9:0] funct,     // {funct7, funct3}
    output wire [3:0] alu_control 
);


endmodule