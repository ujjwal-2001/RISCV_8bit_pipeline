module Control
(
    input wire [6:0] opcode,
    output wire branch,
    output wire mem_read,
    output wire mem_to_reg,
    output wire [1:0] alu_op,
    output wire mem_write,
    output wire alu_src,
    output wire reg_write
);

        

endmodule