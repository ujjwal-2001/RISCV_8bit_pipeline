module ALU 
(
    input wire [7:0] data1,
    input wire [7:0] data2,
    input wire [3:0] ALU_control,
    output wire [7:0] ALU_result,
    output wire zero
);



endmodule